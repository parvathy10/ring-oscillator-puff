`timescale 1ns / 1ps
module top(input [7:0] sel1,input[7:0] sel2,
           input enable,reset,
          output m1out,m2out,
           output [127:0]count_1 , output [127:0]count_2, 
			 output count
          );
  //  wire w1, w2, w3, w4, w5, w6, w7, w8;
       // wire[15:0] w11, w12;
  wire [127:0] din1, din2;
    // wire [7:0] count1; wire [7:0]count2;
 ro1 ro1(enable,din1[0]);
ro2 ro2(enable,din1[1]);
ro3 ro3(enable,din1[2]);
ro4 ro4(enable,din1[3]);
ro5 ro5(enable,din1[4]);
ro6 ro6(enable,din1[5]);
ro7 ro7(enable,din1[6]);
ro8 ro8(enable,din1[7]);
ro9 ro9(enable,din1[8]);
ro10 ro10(enable,din1[9]);
ro11 ro11(enable,din1[10]);
ro12 ro12(enable,din1[11]);
ro13 ro13(enable,din1[12]);
ro14 ro14(enable,din1[13]);
ro15 ro15(enable,din1[14]);
ro16 ro16(enable,din1[15]);
ro17 ro17(enable,din1[16]);
ro18 ro18(enable,din1[17]);
ro19 ro19(enable,din1[18]);
ro20 ro20(enable,din1[19]);
ro21 ro21(enable,din1[20]);
ro22 ro22(enable,din1[21]);
ro23 ro23(enable,din1[22]);
ro24 ro24(enable,din1[23]);
ro25 ro25(enable,din1[24]);
ro26 ro26(enable,din1[25]);
ro27 ro27(enable,din1[26]);
ro28 ro28(enable,din1[27]);
ro29 ro29(enable,din1[28]);
ro30 ro30(enable,din1[29]);
ro31 ro31(enable,din1[30]);
ro32 ro32(enable,din1[31]);
ro33 ro33(enable,din1[32]);
ro34 ro34(enable,din1[33]);
ro35 ro35(enable,din1[34]);
ro36 ro36(enable,din1[35]);
ro37 ro37(enable,din1[36]);
ro38 ro38(enable,din1[37]);
ro39 ro39(enable,din1[38]);
ro40 ro40(enable,din1[39]);
ro41 ro41(enable,din1[40]);
ro42 ro42(enable,din1[41]);
ro43 ro43(enable,din1[42]);
ro44 ro44(enable,din1[43]);
ro45 ro45(enable,din1[44]);
ro46 ro46(enable,din1[45]);
ro47 ro47(enable,din1[46]);
ro48 ro48(enable,din1[47]);
ro49 ro49(enable,din1[48]);
ro50 ro50(enable,din1[49]);
ro51 ro51(enable,din1[50]);
ro52 ro52(enable,din1[51]);
ro53 ro53(enable,din1[52]);
ro54 ro54(enable,din1[53]);
ro55 ro55(enable,din1[54]);
ro56 ro56(enable,din1[55]);
ro57 ro57(enable,din1[56]);
ro58 ro58(enable,din1[57]);
ro59 ro59(enable,din1[58]);
ro60 ro60(enable,din1[59]);
ro61 ro61(enable,din1[60]);
ro62 ro62(enable,din1[61]);
ro63 ro63(enable,din1[62]);
ro64 ro64(enable,din1[63]);
ro65 ro65(enable,din1[64]);
ro66 ro66(enable,din1[65]);
ro67 ro67(enable,din1[66]);
ro68 ro68(enable,din1[67]);
ro69 ro69(enable,din1[68]);
ro70 ro70(enable,din1[69]);
ro71 ro71(enable,din1[70]);
ro72 ro72(enable,din1[71]);
ro73 ro73(enable,din1[72]);
ro74 ro74(enable,din1[73]);
ro75 ro75(enable,din1[74]);
ro76 ro76(enable,din1[75]);
ro77 ro77(enable,din1[76]);
ro78 ro78(enable,din1[77]);
ro79 ro79(enable,din1[78]);
ro80 ro80(enable,din1[79]);
ro81 ro81(enable,din1[80]);
ro82 ro82(enable,din1[81]);
ro83 ro83(enable,din1[82]);
ro84 ro84(enable,din1[83]);
ro85 ro85(enable,din1[84]);
ro86 ro86(enable,din1[85]);
ro87 ro87(enable,din1[86]);
ro88 ro88(enable,din1[87]);
ro89 ro89(enable,din1[88]);
ro90 ro90(enable,din1[89]);
ro91 ro91(enable,din1[90]);
ro92 ro92(enable,din1[91]);
ro93 ro93(enable,din1[92]);
ro94 ro94(enable,din1[93]);
ro95 ro95(enable,din1[94]);
ro96 ro96(enable,din1[95]);
ro97 ro97(enable,din1[96]);
ro98 ro98(enable,din1[97]);
ro99 ro99(enable,din1[98]);
ro100 ro100(enable,din1[99]);
ro101 ro101(enable,din1[100]);
ro102 ro102(enable,din1[101]);
ro103 ro103(enable,din1[102]);
ro104 ro104(enable,din1[103]);
ro105 ro105(enable,din1[104]);
ro106 ro106(enable,din1[105]);
ro107 ro107(enable,din1[106]);
ro108 ro108(enable,din1[107]);
ro109 ro109(enable,din1[108]);
ro110 ro110(enable,din1[109]);
ro111 ro111(enable,din1[110]);
ro112 ro112(enable,din1[111]);
ro113 ro113(enable,din1[112]);
ro114 ro114(enable,din1[113]);
ro115 ro115(enable,din1[114]);
ro116 ro116(enable,din1[115]);
ro117 ro117(enable,din1[116]);
ro118 ro118(enable,din1[117]);
ro119 ro119(enable,din1[118]);
ro120 ro120(enable,din1[119]);
ro121 ro121(enable,din1[120]);
ro122 ro122(enable,din1[121]);
ro123 ro123(enable,din1[122]);
ro124 ro124(enable,din1[123]);
ro125 ro125(enable,din1[124]);
ro126 ro126(enable,din1[125]);
ro127 ro127(enable,din1[126]);
ro128 ro128(enable,din1[127]);



ro1 ro129(enable,din2[0]);
ro2 ro130(enable,din2[1]);
ro3 ro131(enable,din2[2]);
ro4 ro132(enable,din2[3]);
ro5 ro133(enable,din2[4]);
ro6 ro134(enable,din2[5]);
ro7 ro135(enable,din2[6]);
ro8 ro136(enable,din2[7]);
ro9 ro137(enable,din2[8]);
ro10 ro138(enable,din2[9]);
ro11 ro139(enable,din2[10]);
ro12 ro140(enable,din2[11]);
ro13 ro141(enable,din2[12]);
ro14 ro142(enable,din2[13]);
ro15 ro143(enable,din2[14]);
ro16 ro144(enable,din2[15]);
ro17 ro145(enable,din2[16]);
ro18 ro146(enable,din2[17]);
ro19 ro147(enable,din2[18]);
ro20 ro148(enable,din2[19]);
ro21 ro149(enable,din2[20]);
ro22 ro150(enable,din2[21]);
ro23 ro151(enable,din2[22]);
ro24 ro152(enable,din2[23]);
ro25 ro153(enable,din2[24]);
ro26 ro154(enable,din2[25]);
ro27 ro155(enable,din2[26]);
ro28 ro156(enable,din2[27]);
ro29 ro157(enable,din2[28]);
ro30 ro158(enable,din2[29]);
ro31 ro159(enable,din2[30]);
ro32 ro160(enable,din2[31]);
ro33 ro161(enable,din2[32]);
ro34 ro162(enable,din2[33]);
ro35 ro163(enable,din2[34]);
ro36 ro164(enable,din2[35]);
ro37 ro165(enable,din2[36]);
ro38 ro166(enable,din2[37]);
ro39 ro167(enable,din2[38]);
ro40 ro168(enable,din2[39]);
ro41 ro169(enable,din2[40]);
ro42 ro170(enable,din2[41]);
ro43 ro171(enable,din2[42]);
ro44 ro172(enable,din2[43]);
ro45 ro173(enable,din2[44]);
ro46 ro174(enable,din2[45]);
ro47 ro175(enable,din2[46]);
ro48 ro176(enable,din2[47]);
ro49 ro177(enable,din2[48]);
ro50 ro178(enable,din2[49]);
ro51 ro179(enable,din2[50]);
ro52 ro180(enable,din2[51]);
ro53 ro181(enable,din2[52]);
ro54 ro182(enable,din2[53]);
ro55 ro183(enable,din2[54]);
ro56 ro184(enable,din2[55]);
ro57 ro185(enable,din2[56]);
ro58 ro186(enable,din2[57]);
ro59 ro187(enable,din2[58]);
ro60 ro188(enable,din2[59]);
ro61 ro189(enable,din2[60]);
ro62 ro190(enable,din2[61]);
ro63 ro191(enable,din2[62]);
ro64 ro192(enable,din2[63]);
ro65 ro193(enable,din2[64]);
ro66 ro194(enable,din2[65]);
ro67 ro195(enable,din2[66]);
ro68 ro196(enable,din2[67]);
ro69 ro197(enable,din2[68]);
ro70 ro198(enable,din2[69]);
ro71 ro199(enable,din2[70]);
ro72 ro200(enable,din2[71]);
ro73 ro201(enable,din2[72]);
ro74 ro202(enable,din2[73]);
ro75 ro203(enable,din2[74]);
ro76 ro204(enable,din2[75]);
ro77 ro205(enable,din2[76]);
ro78 ro206(enable,din2[77]);
ro79 ro207(enable,din2[78]);
ro80 ro208(enable,din2[79]);
ro81 ro209(enable,din2[80]);
ro82 ro210(enable,din2[81]);
ro83 ro211(enable,din2[82]);
ro84 ro212(enable,din2[83]);
ro85 ro213(enable,din2[84]);
ro86 ro214(enable,din2[85]);
ro87 ro215(enable,din2[86]);
ro88 ro216(enable,din2[87]);
ro89 ro217(enable,din2[88]);
ro90 ro218(enable,din2[89]);
ro91 ro219(enable,din2[90]);
ro92 ro220(enable,din2[91]);
ro93 ro221(enable,din2[92]);
ro94 ro222(enable,din2[93]);
ro95 ro223(enable,din2[94]);
ro96 ro224(enable,din2[95]);
ro97 ro225(enable,din2[96]);
ro98 ro226(enable,din2[97]);
ro99 ro227(enable,din2[98]);
ro100 ro228(enable,din2[99]);
ro101 ro229(enable,din2[100]);
ro102 ro230(enable,din2[101]);
ro103 ro231(enable,din2[102]);
ro104 ro232(enable,din2[103]);
ro105 ro233(enable,din2[104]);
ro106 ro234(enable,din2[105]);
ro107 ro235(enable,din2[106]);
ro108 ro236(enable,din2[107]);
ro109 ro237(enable,din2[108]);
ro110 ro238(enable,din2[109]);
ro111 ro239(enable,din2[110]);
ro112 ro240(enable,din2[111]);
ro113 ro241(enable,din2[112]);
ro114 ro242(enable,din2[113]);
ro115 ro243(enable,din2[114]);
ro116 ro244(enable,din2[115]);
ro117 ro245(enable,din2[116]);
ro118 ro246(enable,din2[117]);
ro119 ro247(enable,din2[118]);
ro120 ro248(enable,din2[119]);
ro121 ro249(enable,din2[120]);
ro122 ro250(enable,din2[121]);
ro123 ro251(enable,din2[122]);
ro124 ro252(enable,din2[123]);
ro125 ro253(enable,din2[124]);
ro126 ro254(enable,din2[125]);
ro127 ro255(enable,din2[126]);
ro128 ro256(enable,din2[127]);
  


   
      mux_16 M1(din1,m1out,sel1 );
      mux_16 M2(din2,m2out ,sel2);
		 
         
				 
         //cac cac(m1out,m2out,enable,reset, count_1, count_2);
			cac2 cac2(m2out,m1out,enable,reset, count_2, count_1);

        comp comp(count_2,count_1,count) ;
			  
            
endmodule
