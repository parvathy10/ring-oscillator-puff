`timescale 1ns/1ps
module ro1(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        nand #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
       
		
endmodule

module ro2(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #2(w1, en, out);
        not #2(w2, w1);
        not #2(w3, w2);
        not #2(w4,w3);
        not #2(w5, w4);
        not #2(out, w5);
        
		
endmodule

module ro3(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;
		
		  
        nand #3(w1, en, out);
        not #3(w2, w1);
        not #3(w3, w2);
        not #3(w4,w3);
        not #3(w5, w4);
        not #3(out, w5);
        
		
endmodule

module ro4(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;
		
		  
        nand #4(w1, en, out);
        not #4(w2, w1);
        not #4(w3, w2);
        not #4(w4,w3);
        not #4(w5, w4);
        not #4(out, w5);
        
		
endmodule

module ro5(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #5(w1, en, out);
        not #5(w2, w1);
        not #5(w3, w2);
        not #5(w4,w3);
        not #5(w5, w4);
        not #5(out, w5);
       
		
endmodule

module ro6(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;
		
		  
        nand #6(w1, en, out);
        not #6(w2, w1);
        not #6(w3, w2);
        not #6(w4,w3);
        not #6(w5, w4);
        not #6(out, w5);
        
endmodule

module ro7(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        nand #7(w1, en, out);
        not #7(w2, w1);
        not #7(w3, w2);
        not #7(w4,w3);
        not #7(w5, w4);
        not #7(out, w5);
       
		
endmodule

module ro8(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #8(w1, en, out);
        not #8(w2, w1);
        not #8(w3, w2);
        not #8(w4,w3);
        not #8(w5, w4);
        not #8(out, w5);
        
		
endmodule
module ro9(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #9(w1, en, out);
        not #9(w2, w1);
        not #9(w3, w2);
        not #9(w4,w3);
        not #9(w5, w4);
        not #9(out, w5);
        
		
endmodule

module ro10(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #10(w1, en, out);
        not #10(w2, w1);
        not #10(w3, w2);
        not #10(w4,w3);
        not #10(w5, w4);
        not #10(out, w5);
        
		
endmodule

module ro11(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #11(w1, en, out);
        not #11(w2, w1);
        not #11(w3, w2);
        not #11(w4,w3);
        not #11(w5, w4);
        not #11(out, w5);
        
		
endmodule

module ro12(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #12(w1, en, out);
        not #12(w2, w1);
        not #12(w3, w2);
        not #12(w4,w3);
        not #12(w5, w4);
        not #12(out, w5);
        
		
endmodule

module ro13(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #13(w1, en, out);
        not #13(w2, w1);
        not #13(w3, w2);
        not #13(w4,w3);
        not #13(w5, w4);
        not #13(out, w5);
        
		
endmodule

module ro14(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #14(w1, en, out);
        not #14(w2, w1);
        not #14(w3, w2);
        not #14(w4,w3);
        not #14(w5, w4);
        not #14(out, w5);
        
		
endmodule

module ro15(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #15(w1, en, out);
        not #15(w2, w1);
        not #15(w3, w2);
        not #15(w4,w3);
        not #15(w5, w4);
        not #15(out, w5);
        
		
endmodule

module ro16(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #16(w1, en, out);
        not #16(w2, w1);
        not #16(w3, w2);
        not #16(w4,w3);
        not #16(w5, w4);
        not #16(out, w5);
        
		
endmodule

module ro17(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #17(w1, en, out);
        not #17(w2, w1);
        not #17(w3, w2);
        not #17(w4,w3);
        not #17(w5, w4);
        not #17(out, w5);
        
		
endmodule

module ro18(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #18(w1, en, out);
        not #18(w2, w1);
        not #18(w3, w2);
        not #18(w4,w3);
        not #18(w5, w4);
        not #18(out, w5);
        
		
endmodule

module ro19(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #19(w1, en, out);
        not #19(w2, w1);
        not #19(w3, w2);
        not #19(w4,w3);
        not #19(w5, w4);
        not #19(out, w5);
        
		
endmodule
  
module ro20(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #20(w1, en, out);
        not #20(w2, w1);
        not #20(w3, w2);
        not #20(w4,w3);
        not #20(w5, w4);
        not #20(out, w5);
        
		
endmodule
  
module ro21(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #21(w1, en, out);
        not #21(w2, w1);
        not #21(w3, w2);
        not #21(w4,w3);
        not #21(w5, w4);
        not #21(out, w5);
        
		
endmodule
  
module ro22(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #22(w1, en, out);
        not #22(w2, w1);
        not #22(w3, w2);
        not #22(w4,w3);
        not #22(w5, w4);
        not #22(out, w5);
        
		
endmodule
  
module ro23(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #23(w1, en, out);
        not #23(w2, w1);
        not #23(w3, w2);
        not #23(w4,w3);
        not #23(w5, w4);
        not #23(out, w5);
        
		
endmodule
  
module ro24(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #24(w1, en, out);
        not #24(w2, w1);
        not #24(w3, w2);
        not #24(w4,w3);
        not #24(w5, w4);
        not #24(out, w5);
        
		
endmodule
  
module ro25(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #25(w1, en, out);
        not #25(w2, w1);
        not #25(w3, w2);
        not #25(w4,w3);
        not #25(w5, w4);
        not #25(out, w5);
        
		
endmodule
  
module ro26(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #26(w1, en, out);
        not #26(w2, w1);
        not #26(w3, w2);
        not #26(w4,w3);
        not #26(w5, w4);
        not #26(out, w5);
        
		
endmodule
  
module ro27(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #27(w1, en, out);
        not #27(w2, w1);
        not #27(w3, w2);
        not #27(w4,w3);
        not #27(w5, w4);
        not #27(out, w5);
        
		
endmodule
  
module ro28(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #28(w1, en, out);
        not #28(w2, w1);
        not #28(w3, w2);
        not #28(w4,w3);
        not #28(w5, w4);
        not #28(out, w5);
        
		
endmodule
  
module ro29(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #29(w1, en, out);
        not #29(w2, w1);
        not #29(w3, w2);
        not #29(w4,w3);
        not #29(w5, w4);
        not #29(out, w5);
        
		
endmodule
  
module ro30(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #30(w1, en, out);
        not #30(w2, w1);
        not #30(w3, w2);
        not #30(w4,w3);
        not #30(w5, w4);
        not #30(out, w5);
        
		
endmodule
  
module ro31(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #31(w1, en, out);
        not #31(w2, w1);
        not #31(w3, w2);
        not #31(w4,w3);
        not #31(w5, w4);
        not #31(out, w5);
        
		
endmodule
  
module ro32(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #32(w1, en, out);
        not #32(w2, w1);
        not #32(w3, w2);
        not #32(w4,w3);
        not #32(w5, w4);
        not #32(out, w5);
        
		
endmodule
  
module ro33(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #33(w1, en, out);
        not #33(w2, w1);
        not #33(w3, w2);
        not #33(w4,w3);
        not #33(w5, w4);
        not #33(out, w5);
        
		
endmodule
  
module ro34(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #34(w1, en, out);
        not #34(w2, w1);
        not #34(w3, w2);
        not #34(w4,w3);
        not #34(w5, w4);
        not #34(out, w5);
        
		
endmodule
  
module ro35(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #35(w1, en, out);
        not #35(w2, w1);
        not #35(w3, w2);
        not #35(w4,w3);
        not #35(w5, w4);
        not #35(out, w5);
        
		
endmodule
  
module ro36(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #36(w1, en, out);
        not #36(w2, w1);
        not #36(w3, w2);
        not #36(w4,w3);
        not #36(w5, w4);
        not #36(out, w5);
        
		
endmodule
  
module ro37(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #37(w1, en, out);
        not #37(w2, w1);
        not #37(w3, w2);
        not #37(w4,w3);
        not #37(w5, w4);
        not #37(out, w5);
        
		
endmodule
  
module ro38(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #38(w1, en, out);
        not #38(w2, w1);
        not #38(w3, w2);
        not #38(w4,w3);
        not #38(w5, w4);
        not #38(out, w5);
        
		
endmodule
  
module ro39(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #39(w1, en, out);
        not #39(w2, w1);
        not #39(w3, w2);
        not #39(w4,w3);
        not #39(w5, w4);
        not #39(out, w5);
        
		
endmodule
  
module ro40(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #40(w1, en, out);
        not #40(w2, w1);
        not #40(w3, w2);
        not #40(w4,w3);
        not #40(w5, w4);
        not #40(out, w5);
        
		
endmodule
  
module ro41(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #41(w1, en, out);
        not #41(w2, w1);
        not #41(w3, w2);
        not #41(w4,w3);
        not #41(w5, w4);
        not #41(out, w5);
        
		
endmodule
  
module ro42(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #42(w1, en, out);
        not #42(w2, w1);
        not #42(w3, w2);
        not #42(w4,w3);
        not #42(w5, w4);
        not #42(out, w5);
        
		
endmodule
  
module ro43(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #43(w1, en, out);
        not #43(w2, w1);
        not #43(w3, w2);
        not #43(w4,w3);
        not #43(w5, w4);
        not #43(out, w5);
        
		
endmodule
  
module ro44(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #44(w1, en, out);
        not #44(w2, w1);
        not #44(w3, w2);
        not #44(w4,w3);
        not #44(w5, w4);
        not #44(out, w5);
        
		
endmodule
  
module ro45(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #45(w1, en, out);
        not #45(w2, w1);
        not #45(w3, w2);
        not #45(w4,w3);
        not #45(w5, w4);
        not #45(out, w5);
        
		
endmodule
  
module ro46(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #46(w1, en, out);
        not #46(w2, w1);
        not #46(w3, w2);
        not #46(w4,w3);
        not #46(w5, w4);
        not #46(out, w5);
        
		
endmodule
  
module ro47(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #47(w1, en, out);
        not #47(w2, w1);
        not #47(w3, w2);
        not #47(w4,w3);
        not #47(w5, w4);
        not #47(out, w5);
        
		
endmodule
  
module ro48(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #48(w1, en, out);
        not #48(w2, w1);
        not #48(w3, w2);
        not #48(w4,w3);
        not #48(w5, w4);
        not #48(out, w5);
        
		
endmodule
  
module ro49(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #49(w1, en, out);
        not #49(w2, w1);
        not #49(w3, w2);
        not #49(w4,w3);
        not #49(w5, w4);
        not #49(out, w5);
        
		
endmodule
  
module ro50(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #50(w1, en, out);
        not #50(w2, w1);
        not #50(w3, w2);
        not #50(w4,w3);
        not #50(w5, w4);
        not #50(out, w5);
        
		
endmodule
  
module ro51(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #51(w1, en, out);
        not #51(w2, w1);
        not #51(w3, w2);
        not #51(w4,w3);
        not #51(w5, w4);
        not #51(out, w5);
        
		
endmodule
  
module ro52(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #52(w1, en, out);
        not #52(w2, w1);
        not #52(w3, w2);
        not #52(w4,w3);
        not #52(w5, w4);
        not #52(out, w5);
        
		
endmodule
  
module ro53(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #53(w1, en, out);
        not #53(w2, w1);
        not #53(w3, w2);
        not #53(w4,w3);
        not #53(w5, w4);
        not #53(out, w5);
        
		
endmodule
  
module ro54(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #54(w1, en, out);
        not #54(w2, w1);
        not #54(w3, w2);
        not #54(w4,w3);
        not #54(w5, w4);
        not #54(out, w5);
        
		
endmodule
  
module ro55(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #55(w1, en, out);
        not #55(w2, w1);
        not #55(w3, w2);
        not #55(w4,w3);
        not #55(w5, w4);
        not #55(out, w5);
        
		
endmodule
  
module ro56(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #56(w1, en, out);
        not #56(w2, w1);
        not #56(w3, w2);
        not #56(w4,w3);
        not #56(w5, w4);
        not #56(out, w5);
        
		
endmodule
  
module ro57(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #57(w1, en, out);
        not #57(w2, w1);
        not #57(w3, w2);
        not #57(w4,w3);
        not #57(w5, w4);
        not #57(out, w5);
        
		
endmodule
  
module ro58(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #58(w1, en, out);
        not #58(w2, w1);
        not #58(w3, w2);
        not #58(w4,w3);
        not #58(w5, w4);
        not #58(out, w5);
        
		
endmodule
  
module ro59(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #59(w1, en, out);
        not #59(w2, w1);
        not #59(w3, w2);
        not #59(w4,w3);
        not #59(w5, w4);
        not #59(out, w5);
        
		
endmodule
  
module ro60(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #60(w1, en, out);
        not #60(w2, w1);
        not #60(w3, w2);
        not #60(w4,w3);
        not #60(w5, w4);
        not #60(out, w5);
        
		
endmodule
  
module ro61(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #61(w1, en, out);
        not #61(w2, w1);
        not #61(w3, w2);
        not #61(w4,w3);
        not #61(w5, w4);
        not #61(out, w5);
        
		
endmodule
  
module ro62(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #62(w1, en, out);
        not #62(w2, w1);
        not #62(w3, w2);
        not #62(w4,w3);
        not #62(w5, w4);
        not #62(out, w5);
        
		
endmodule
  
module ro63(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #63(w1, en, out);
        not #63(w2, w1);
        not #63(w3, w2);
        not #63(w4,w3);
        not #63(w5, w4);
        not #63(out, w5);
        
		
endmodule
  
module ro64(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #64(w1, en, out);
        not #64(w2, w1);
        not #64(w3, w2);
        not #64(w4,w3);
        not #64(w5, w4);
        not #64(out, w5);
        
		
endmodule
  
module ro65(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #65(w1, en, out);
        not #65(w2, w1);
        not #65(w3, w2);
        not #65(w4,w3);
        not #65(w5, w4);
        not #65(out, w5);
        
		
endmodule
  
module ro66(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #66(w1, en, out);
        not #66(w2, w1);
        not #66(w3, w2);
        not #66(w4,w3);
        not #66(w5, w4);
        not #66(out, w5);
        
		
endmodule
  
module ro67(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #67(w1, en, out);
        not #67(w2, w1);
        not #67(w3, w2);
        not #67(w4,w3);
        not #67(w5, w4);
        not #67(out, w5);
        
		
endmodule
  
module ro68(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #68(w1, en, out);
        not #68(w2, w1);
        not #68(w3, w2);
        not #68(w4,w3);
        not #68(w5, w4);
        not #68(out, w5);
        
		
endmodule
  
module ro69(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #69(w1, en, out);
        not #69(w2, w1);
        not #69(w3, w2);
        not #69(w4,w3);
        not #69(w5, w4);
        not #69(out, w5);
        
		
endmodule
  
module ro70(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #70(w1, en, out);
        not #70(w2, w1);
        not #70(w3, w2);
        not #70(w4,w3);
        not #70(w5, w4);
        not #70(out, w5);
        
		
endmodule
  
module ro71(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #71(w1, en, out);
        not #71(w2, w1);
        not #71(w3, w2);
        not #71(w4,w3);
        not #71(w5, w4);
        not #71(out, w5);
        
		
endmodule
  
module ro72(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #72(w1, en, out);
        not #72(w2, w1);
        not #72(w3, w2);
        not #72(w4,w3);
        not #72(w5, w4);
        not #72(out, w5);
        
		
endmodule
  
module ro73(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #73(w1, en, out);
        not #73(w2, w1);
        not #73(w3, w2);
        not #73(w4,w3);
        not #73(w5, w4);
        not #73(out, w5);
        
		
endmodule
  
module ro74(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #74(w1, en, out);
        not #74(w2, w1);
        not #74(w3, w2);
        not #74(w4,w3);
        not #74(w5, w4);
        not #74(out, w5);
        
		
endmodule
  
module ro75(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #75(w1, en, out);
        not #75(w2, w1);
        not #75(w3, w2);
        not #75(w4,w3);
        not #75(w5, w4);
        not #75(out, w5);
        
		
endmodule
  
module ro76(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #76(w1, en, out);
        not #76(w2, w1);
        not #76(w3, w2);
        not #76(w4,w3);
        not #76(w5, w4);
        not #76(out, w5);
        
		
endmodule
  
module ro77(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #77(w1, en, out);
        not #77(w2, w1);
        not #77(w3, w2);
        not #77(w4,w3);
        not #77(w5, w4);
        not #77(out, w5);
        
		
endmodule
  
module ro78(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #78(w1, en, out);
        not #78(w2, w1);
        not #78(w3, w2);
        not #78(w4,w3);
        not #78(w5, w4);
        not #78(out, w5);
        
		
endmodule
  
module ro79(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #79(w1, en, out);
        not #79(w2, w1);
        not #79(w3, w2);
        not #79(w4,w3);
        not #79(w5, w4);
        not #79(out, w5);
        
		
endmodule
  
module ro80(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #80(w1, en, out);
        not #80(w2, w1);
        not #80(w3, w2);
        not #80(w4,w3);
        not #80(w5, w4);
        not #80(out, w5);
        
		
endmodule
  
module ro81(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #81(w1, en, out);
        not #81(w2, w1);
        not #81(w3, w2);
        not #81(w4,w3);
        not #81(w5, w4);
        not #81(out, w5);
        
		
endmodule
  
module ro82(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #82(w1, en, out);
        not #82(w2, w1);
        not #82(w3, w2);
        not #82(w4,w3);
        not #82(w5, w4);
        not #82(out, w5);
        
		
endmodule
  
module ro83(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #83(w1, en, out);
        not #83(w2, w1);
        not #83(w3, w2);
        not #83(w4,w3);
        not #83(w5, w4);
        not #83(out, w5);
        
		
endmodule
  
module ro84(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #84(w1, en, out);
        not #84(w2, w1);
        not #84(w3, w2);
        not #84(w4,w3);
        not #84(w5, w4);
        not #84(out, w5);
        
		
endmodule
  
module ro85(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #85(w1, en, out);
        not #85(w2, w1);
        not #85(w3, w2);
        not #85(w4,w3);
        not #85(w5, w4);
        not #85(out, w5);
        
		
endmodule
  
module ro86(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #86(w1, en, out);
        not #86(w2, w1);
        not #86(w3, w2);
        not #86(w4,w3);
        not #86(w5, w4);
        not #86(out, w5);
        
		
endmodule
  
module ro87(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #87(w1, en, out);
        not #87(w2, w1);
        not #87(w3, w2);
        not #87(w4,w3);
        not #87(w5, w4);
        not #87(out, w5);
        
		
endmodule
  
module ro88(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #88(w1, en, out);
        not #88(w2, w1);
        not #88(w3, w2);
        not #88(w4,w3);
        not #88(w5, w4);
        not #88(out, w5);
        
		
endmodule
  
module ro89(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #89(w1, en, out);
        not #89(w2, w1);
        not #89(w3, w2);
        not #89(w4,w3);
        not #89(w5, w4);
        not #89(out, w5);
        
		
endmodule
  
module ro90(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #90(w1, en, out);
        not #90(w2, w1);
        not #90(w3, w2);
        not #90(w4,w3);
        not #90(w5, w4);
        not #90(out, w5);
        
		
endmodule
  
module ro91(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #91(w1, en, out);
        not #91(w2, w1);
        not #91(w3, w2);
        not #91(w4,w3);
        not #91(w5, w4);
        not #91(out, w5);
        
		
endmodule
  
module ro92(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #92(w1, en, out);
        not #92(w2, w1);
        not #92(w3, w2);
        not #92(w4,w3);
        not #92(w5, w4);
        not #92(out, w5);
        
		
endmodule
  
module ro93(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #93(w1, en, out);
        not #93(w2, w1);
        not #93(w3, w2);
        not #93(w4,w3);
        not #93(w5, w4);
        not #93(out, w5);
        
		
endmodule
  
module ro94(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #94(w1, en, out);
        not #94(w2, w1);
        not #94(w3, w2);
        not #94(w4,w3);
        not #94(w5, w4);
        not #94(out, w5);
        
		
endmodule
  
module ro95(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #95(w1, en, out);
        not #95(w2, w1);
        not #95(w3, w2);
        not #95(w4,w3);
        not #95(w5, w4);
        not #95(out, w5);
        
		
endmodule
  
module ro96(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #96(w1, en, out);
        not #96(w2, w1);
        not #96(w3, w2);
        not #96(w4,w3);
        not #96(w5, w4);
        not #96(out, w5);
        
		
endmodule
  
module ro97(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #97(w1, en, out);
        not #97(w2, w1);
        not #97(w3, w2);
        not #97(w4,w3);
        not #97(w5, w4);
        not #97(out, w5);
        
		
endmodule
  
module ro98(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #98(w1, en, out);
        not #98(w2, w1);
        not #98(w3, w2);
        not #98(w4,w3);
        not #98(w5, w4);
        not #98(out, w5);
        
		
endmodule
  
module ro99(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #99(w1, en, out);
        not #99(w2, w1);
        not #99(w3, w2);
        not #99(w4,w3);
        not #99(w5, w4);
        not #99(out, w5);
        
		
endmodule
  
module ro100(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #100(w1, en, out);
        not #100(w2, w1);
        not #100(w3, w2);
        not #100(w4,w3);
        not #100(w5, w4);
        not #100(out, w5);
        
		
endmodule
  
module ro101(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #101(w1, en, out);
        not #101(w2, w1);
        not #101(w3, w2);
        not #101(w4,w3);
        not #101(w5, w4);
        not #101(out, w5);
        
		
endmodule
  
module ro102(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #102(w1, en, out);
        not #102(w2, w1);
        not #102(w3, w2);
        not #102(w4,w3);
        not #102(w5, w4);
        not #102(out, w5);
        
		
endmodule
  
module ro103(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #103(w1, en, out);
        not #103(w2, w1);
        not #103(w3, w2);
        not #103(w4,w3);
        not #103(w5, w4);
        not #103(out, w5);
        
		
endmodule
  
module ro104(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #104(w1, en, out);
        not #104(w2, w1);
        not #104(w3, w2);
        not #104(w4,w3);
        not #104(w5, w4);
        not #104(out, w5);
        
		
endmodule
  
module ro105(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #105(w1, en, out);
        not #105(w2, w1);
        not #105(w3, w2);
        not #105(w4,w3);
        not #105(w5, w4);
        not #105(out, w5);
        
		
endmodule
  
module ro106(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #106(w1, en, out);
        not #106(w2, w1);
        not #106(w3, w2);
        not #106(w4,w3);
        not #106(w5, w4);
        not #106(out, w5);
        
		
endmodule
  
module ro107(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #107(w1, en, out);
        not #107(w2, w1);
        not #107(w3, w2);
        not #107(w4,w3);
        not #107(w5, w4);
        not #107(out, w5);
        
		
endmodule
  
module ro108(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #108(w1, en, out);
        not #108(w2, w1);
        not #108(w3, w2);
        not #108(w4,w3);
        not #108(w5, w4);
        not #108(out, w5);
        
		
endmodule
  
module ro109(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #109(w1, en, out);
        not #109(w2, w1);
        not #109(w3, w2);
        not #109(w4,w3);
        not #109(w5, w4);
        not #109(out, w5);
        
		
endmodule
  
  
module ro110(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #110(w1, en, out);
        not #110(w2, w1);
        not #110(w3, w2);
        not #110(w4,w3);
        not #110(w5, w4);
        not #110(out, w5);
        
		
endmodule
  
  
module ro111(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #111(w1, en, out);
        not #111(w2, w1);
        not #111(w3, w2);
        not #111(w4,w3);
        not #111(w5, w4);
        not #111(out, w5);
        
		
endmodule
  
module ro112(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #112(w1, en, out);
        not #112(w2, w1);
        not #112(w3, w2);
        not #112(w4,w3);
        not #112(w5, w4);
        not #112(out, w5);
        
		
endmodule
  
module ro113(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #113(w1, en, out);
        not #113(w2, w1);
        not #113(w3, w2);
        not #113(w4,w3);
        not #113(w5, w4);
        not #113(out, w5);
        
		
endmodule
  
module ro114(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #114(w1, en, out);
        not #114(w2, w1);
        not #114(w3, w2);
        not #114(w4,w3);
        not #114(w5, w4);
        not #114(out, w5);
        
		
endmodule
  
module ro115(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #115(w1, en, out);
        not #115(w2, w1);
        not #115(w3, w2);
        not #115(w4,w3);
        not #115(w5, w4);
        not #115(out, w5);
        
		
endmodule
  
module ro116(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #116(w1, en, out);
        not #116(w2, w1);
        not #116(w3, w2);
        not #116(w4,w3);
        not #116(w5, w4);
        not #116(out, w5);
        
		
endmodule
  
module ro117(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #117(w1, en, out);
        not #117(w2, w1);
        not #117(w3, w2);
        not #117(w4,w3);
        not #117(w5, w4);
        not #117(out, w5);
        
		
endmodule
  
module ro118(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #118(w1, en, out);
        not #118(w2, w1);
        not #118(w3, w2);
        not #118(w4,w3);
        not #118(w5, w4);
        not #118(out, w5);
        
		
endmodule
  
module ro119(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #119(w1, en, out);
        not #119(w2, w1);
        not #119(w3, w2);
        not #119(w4,w3);
        not #119(w5, w4);
        not #119(out, w5);
        
		
endmodule
  
module ro120(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #120(w1, en, out);
        not #120(w2, w1);
        not #120(w3, w2);
        not #120(w4,w3);
        not #120(w5, w4);
        not #120(out, w5);
        
		
endmodule
  
module ro121(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #121(w1, en, out);
        not #121(w2, w1);
        not #121(w3, w2);
        not #121(w4,w3);
        not #121(w5, w4);
        not #121(out, w5);
        
		
endmodule
  
module ro122(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #122(w1, en, out);
        not #122(w2, w1);
        not #122(w3, w2);
        not #122(w4,w3);
        not #122(w5, w4);
        not #122(out, w5);
        
		
endmodule
  
module ro123(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #123(w1, en, out);
        not #123(w2, w1);
        not #123(w3, w2);
        not #123(w4,w3);
        not #123(w5, w4);
        not #123(out, w5);
        
		
endmodule
  
module ro124(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #124(w1, en, out);
        not #124(w2, w1);
        not #124(w3, w2);
        not #124(w4,w3);
        not #124(w5, w4);
        not #124(out, w5);
        
		
endmodule
  
module ro125(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #125(w1, en, out);
        not #125(w2, w1);
        not #125(w3, w2);
        not #125(w4,w3);
        not #125(w5, w4);
        not #125(out, w5);
        
		
endmodule
  
module ro126(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #126(w1, en, out);
        not #126(w2, w1);
        not #126(w3, w2);
        not #126(w4,w3);
        not #126(w5, w4);
        not #126(out, w5);
        
		
endmodule

module ro127(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #127(w1, en, out);
        not #127(w2, w1);
        not #127(w3, w2);
        not #127(w4,w3);
        not #127(w5, w4);
        not #127(out, w5);
        
		
endmodule

module ro128(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5; 
		
		  
        nand #128(w1, en, out);
        not #128(w2, w1);
        not #128(w3, w2);
        not #128(w4,w3);
        not #128(w5, w4);
        not #128(out, w5);
        
		
endmodule




